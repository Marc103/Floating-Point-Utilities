package golden_models_pkg;
    `include "FpModel32.sv"
endpackage
package scoreboards_pkg;
    `include "FpScoreboard32.sv"
endpackage
package monitors_pkg;
    `include "monitors_pkg.sv"
endpackage
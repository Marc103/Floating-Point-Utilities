package monitors_pkg;
    `include "FpMonitor32.sv"
    `include "WindowFetcherMonitor.sv"
endpackage
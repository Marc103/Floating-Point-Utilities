package generators_pkg;
    `include "FpGenerator32.sv"
    `include "ImageGenerator.sv"
    `include "ConvolutionFloatingPointGenerator.sv"
endpackage
package generators_pkg;
    `include "FpGenerator32.sv"
endpackage
package drivers_pkg;
    `include "FpDriver32.sv"
    `include "WindowFetcherDriver.sv"
    `include "ConvolutionFloatingPointDriver.sv"
endpackage
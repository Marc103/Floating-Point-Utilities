package monitors_pkg;
    `include "FpMonitor32.sv"
endpackage
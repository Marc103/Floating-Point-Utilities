package golden_models_pkg;
    `include "FpModel32.sv"
    `include "WindowFetcherModel.sv"
    `include "ConvolutionFloatingPointModel32.sv"
endpackage
package scoreboards_pkg;
    `include "FpScoreboard32.sv"
    `include "WindowFetcherScoreboard.sv"
endpackage
package drivers_pkg;
    `include "FpDriver32.sv"
endpackage
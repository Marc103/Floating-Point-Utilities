package drivers_pkg;
    `include "FpDriver32.sv"
    `include "WindowFetcherDriver.sv"
endpackage
package scoreboards_pkg;
    `include "FpScoreboard32.sv"
    `include "WindowFetcherScoreboard.sv"
    `include "ConvolutionFloatingPointScoreboard32.sv"
endpackage
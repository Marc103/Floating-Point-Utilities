package interfaces_pkg;
    `include "floating_point_inf.svh"
endpackage
package monitors_pkg;
    `include "FpMonitor32.sv"
    `include "WindowFetcherMonitor.sv"
    `include "ConvolutionFloatingPointMonitor.sv"
    `include "DualImageMonitor.sv"
endpackage
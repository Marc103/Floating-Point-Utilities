package FpScoreboard32;
    `include "FpScoreboard32.sv"
endpackage
package utilities_pkg;
    `include "TriggerableQueue.sv"
    `include "TriggerableQueueBroadcaster.sv"
    `include "FloatingPoint.sv"
    `include "Image.sv"
endpackage